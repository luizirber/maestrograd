An�lise CC, Lista 3, Exerc�cio 3
L1 0 2 10mH IC=90mA
R1 2 1 20
C1 1 0 2uF IC=-10V
.TRAN 20u 5000u UIC
.PROBE
.END